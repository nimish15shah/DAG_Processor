
`ifndef CROSSBAR_DEF
  `define CROSSBAR_DEF

`endif //CROSSBAR_DEF
