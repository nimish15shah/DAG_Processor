`include "../proces"
